LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY ov7670_capture IS
    PORT (
	
	    --����� ����� ������
		
        clk : IN STD_LOGIC; --���� ������ ������ (100 ���)
        rst : IN STD_LOGIC;  -- �����
        config_finished : IN STD_LOGIC; --��� ����� "������ ������"
		
		
        -- ����� ������
        --camera signals  
		
        ov7670_vsync : IN STD_LOGIC; -- ����� �����  ,������ ����
        ov7670_href : IN STD_LOGIC; --����� ����,������ �����
        ov7670_pclk : IN STD_LOGIC; --�������� ������ �� ����,���� ��������
        ov7670_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0); --����� ������
		
		--����� ���� ������
		
        start : IN STD_LOGIC;
        frame_finished_o : OUT STD_LOGIC; --��� �����,������ �����
    
        --����� ������� �RAM 
        --frame_buffer signals
		
        wea : OUT STD_LOGIC_VECTOR(0 DOWNTO 0); --����� ����!
        dina : OUT STD_LOGIC_VECTOR(11 DOWNTO 0); -- ������ �����,12 ���
        addra : OUT STD_LOGIC_VECTOR(18 DOWNTO 0) --����� �����
    );
	
END ov7670_capture;

ARCHITECTURE rtl OF ov7670_capture IS
ARCHITECTURE rtl OF ov7670_capture IS
ARCHITECTURE rtl OF ov7670_capture IS

    -- === 1. ����� ������ (State Machine) ===
    TYPE state_type IS (
        idle,                -- ��� �����
        start_capturing,     -- ����� �����
        wait_for_new_frame,  -- ����� ������� ����
        frame_finished,      -- ���� �����
        capture_line,        -- ����� ������ ����
        capture_rgb_byte,    -- ����� ���� ������
        write_to_bram        -- ����� ���� ���� ������
    );

    -- === 2. ������� ������� (Synchronized Signals) ===
    -- �����: ����� ����� ������ �� ������ ����� �� �-FPGA
    -- �� ��� ���� ��� ��� ����-������ (sync1, sync2) ��� ����� ��-������
    
    -- ������ ��� �-VSYNC (����� �����)
    SIGNAL vsync_sync1, vsync_sync2, vsync_prev : STD_LOGIC := '0';
    
    -- ������ ��� �-HREF (����� ����)
    SIGNAL href_sync1, href_sync2, href_prev : STD_LOGIC := '0';
    
    -- ������ ��� �-PCLK (���� �������� - ��� �������� ���� ���� ���� ���)
    SIGNAL pclk_sync1, pclk_sync2, pclk_prev : STD_LOGIC := '0';
    
    -- ������ ����� ����� (Data Bus) - 
    -- �� 8 ������ �� ���� ������ ����� ������ ��� ��� ���� "���" ���� ����
    SIGNAL data_sync1, data_sync2 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');

    -- === 3. ������� ������ ������� (Edge Detection) ===
    -- ����� ����� �-'1' ������ ���� ��� ����� ������ �����
    
    SIGNAL vsync_falling_edge, vsync_rising_edge : STD_LOGIC := '0';
    SIGNAL href_rising_edge, href_falling_edge : STD_LOGIC := '0';
    SIGNAL pclk_rising_edge : STD_LOGIC := '0'; -- ���� ������ ��� ������ �����

    -- === 4. ���� ������� (Registers Record) ===
    TYPE reg_type IS RECORD
        state : state_type;
        href_cnt : INTEGER RANGE 0 TO 500;          -- ���� ����� (�� 480)
        rgb_reg : STD_LOGIC_VECTOR(15 DOWNTO 0);     -- ���� ���� ������ (16 ���)
        pixel_reg : INTEGER RANGE 0 TO 650;         -- ���� ������� ����� (�� 640)
        bram_address : UNSIGNED(18 DOWNTO 0);        -- ����� �������
        line_started : STD_LOGIC;                    -- ���: ��� ������ ����?
    END RECORD reg_type;

	
	-- === 5. ���� ������ (Initialization Constant) -  ===
    -- ��� "�����" �� ���� �������. �������� Reset, ����� ������� �� �� �������.
    CONSTANT INIT_REG_FILE : reg_type := (
        state => idle,                          -- ������� ���� �����
        href_cnt => 0,                          -- ����� ���� �����
        rgb_reg => (OTHERS => '0'),             -- ����� ���� ���� (��� �����)
        pixel_reg => 0,                         -- ����� ���� �������
        bram_address => (OTHERS => '0'),        -- ����� ����� ������� ������ (0)
        line_started => '0'                     -- ����� ��� ����
    );

    -- === 6. ������ ������� (Registers) ===
    -- ��� ����� ������� ����� ������� ����� ��� ����� �� �������� ��� ������
    SIGNAL reg : reg_type := INIT_REG_FILE;      -- ���� ������
    SIGNAL reg_next : reg_type := INIT_REG_FILE; -- ���� ���
	
	
BEGIN

-- === ����� ������ ������� ===
    -- ���� STD_LOGIC_VECTOR ������ ������� (BRAM) ����.
    addra <= STD_LOGIC_VECTOR(reg.bram_address);

    -- === ������ ����� ����� (Edge Detection) ===
    -- ������ �� ��� ������ (Concurrent) ����� ������� ������ ���������.
    -- ��� ����� ��� ���� ������ �������� (sync2) ���� ���� ������ ����� ����� (prev).

    -- ����� ����� VSYNC (�-1 �-0):
    -- ��� ���� ������ ��� ������ ����� ������ ���� ������ ����� (Active Video).
    vsync_falling_edge <= '1' WHEN vsync_prev = '1' AND vsync_sync2 = '0' ELSE '0';

    -- ����� ����� VSYNC (�-0 �-1):
    -- ���� ������� ������� ������� ���� "��" (V-Blank).
    vsync_rising_edge <= '1' WHEN vsync_prev = '0' AND vsync_sync2 = '1' ELSE '0';

    -- ����� ����� HREF (�-0 �-1):
    -- ���� ����� ���� ������ �������� ����� ������� �����.
    href_rising_edge <= '1' WHEN href_prev = '0' AND href_sync2 = '1' ELSE '0';

    -- ����� ����� HREF (�-1 �-0):
    -- ���� ������ �������.
    href_falling_edge <= '1' WHEN href_prev = '1' AND href_sync2 = '0' ELSE '0';

    -- ����� ����� PCLK (�-0 �-1):
    -- ��� "�����" �� �����. ���� ��� ����� ������ ����� ������ ����� �-DATA ��� ���� ����� ������.
    pclk_rising_edge <= '1' WHEN pclk_prev = '0' AND pclk_sync2 = '1' ELSE '0';

    sync : PROCESS (clk, rst)
    BEGIN
        IF rising_edge(clk) THEN
            IF rst = '1' THEN
                reg <= INIT_REG_FILE;
                vsync_sync1 <= '0'; vsync_sync2 <= '0'; vsync_prev <= '0';
                href_sync1 <= '0'; href_sync2 <= '0'; href_prev <= '0';
                pclk_sync1 <= '0'; pclk_sync2 <= '0'; pclk_prev <= '0';
                data_sync1 <= (OTHERS => '0'); data_sync2 <= (OTHERS => '0');
            ELSE
                -- Double buffer for metastability
                vsync_sync1 <= ov7670_vsync; vsync_sync2 <= vsync_sync1; vsync_prev <= vsync_sync2;
                href_sync1 <= ov7670_href;   href_sync2 <= href_sync1;   href_prev <= href_sync2;
                pclk_sync1 <= ov7670_pclk;   pclk_sync2 <= pclk_sync1;   pclk_prev <= pclk_sync2;
                data_sync1 <= ov7670_data;   data_sync2 <= data_sync1;
                
                -- Update registers
                reg <= reg_next;
            END IF;
        END IF;
    END PROCESS;

    comb : PROCESS (reg, data_sync2, pclk_rising_edge, href_rising_edge, href_sync2, start, vsync_falling_edge, vsync_rising_edge, config_finished)
    BEGIN
        reg_next <= reg;
        frame_finished_o <= '0';
        wea <= "0";
        dina <= (OTHERS => '0');
        
        CASE reg.state IS

            WHEN idle =>
                IF start = '1' AND config_finished = '1' THEN
                    reg_next.bram_address <= (OTHERS => '0');
                    reg_next.state <= wait_for_new_frame;
                END IF;

            WHEN wait_for_new_frame =>
                IF vsync_falling_edge = '1' THEN
                    reg_next.href_cnt <= 0;
                    reg_next.bram_address <= (OTHERS => '0'); -- ��� ����� BRAM
                    reg_next.line_started <= '0';
                    reg_next.state <= start_capturing;
                END IF;

            WHEN start_capturing =>
                -- �� �� ����� ����� �� ������ �-HREF ����
                IF href_sync2 = '1' AND reg.line_started = '0' THEN
                    reg_next.pixel_reg <= 0;
					reg_next.bram_address <= to_unsigned(reg.href_cnt * 640, 19);
                    reg_next.line_started <= '1';
                    reg_next.state <= capture_line;
                ELSIF href_sync2 = '0' THEN
                    -- HREF �� ����, ��� �� ����
                    reg_next.line_started <= '0';
                END IF;

            WHEN capture_line =>
                -- ���� �-HREF ����� ���� ��� �� ���� ������
                IF href_sync2 = '1' AND pclk_rising_edge = '1' AND reg.pixel_reg < 640 THEN
                    reg_next.rgb_reg(15 DOWNTO 8) <= data_sync2;
                    reg_next.state <= capture_rgb_byte;
                ELSIF href_sync2 = '0' THEN
                    -- HREF ����, ���� �� �����
                    reg_next.href_cnt <= reg.href_cnt + 1;
                    reg_next.line_started <= '0';
                    IF reg.href_cnt = 479 THEN
                        reg_next.state <= frame_finished;
                    ELSE
                        reg_next.state <= start_capturing;
                    END IF;
                END IF;

            WHEN capture_rgb_byte =>
                IF href_sync2 = '1' AND pclk_rising_edge = '1' AND reg.pixel_reg < 640 THEN
                    reg_next.rgb_reg(7 DOWNTO 0) <= data_sync2;
                    reg_next.pixel_reg <= reg.pixel_reg + 1;
                    reg_next.state <= write_to_bram;
                ELSIF href_sync2 = '0' THEN
                    -- HREF ����, ���� �� �����
                    reg_next.href_cnt <= reg.href_cnt + 1;
                    reg_next.line_started <= '0';
                    IF reg.href_cnt = 479 THEN
                        reg_next.state <= frame_finished;
                    ELSE
                        reg_next.state <= start_capturing;
                    END IF;
                END IF;
                
            WHEN write_to_bram =>
                -- ���� �� �� �� ����� ����
                IF reg.pixel_reg <= 640 AND reg.href_cnt < 480 THEN
                    wea <= "1";
                    dina <= reg.rgb_reg(11 DOWNTO 0);
                    reg_next.bram_address <= reg.bram_address + 1;
                END IF;
                
                -- ���� �� ������ �� �����
                IF reg.pixel_reg >= 640 THEN
                    reg_next.href_cnt <= reg.href_cnt + 1;
                    reg_next.line_started <= '0';
                    IF reg.href_cnt >= 479 THEN
                        reg_next.state <= frame_finished;
                    ELSE
                        reg_next.state <= start_capturing;
                    END IF;
                ELSE
                    reg_next.state <= capture_line;
                END IF;
                
            WHEN frame_finished =>
                frame_finished_o <= '1';
                reg_next.rgb_reg <= (OTHERS => '0');
				reg_next.href_cnt <= 0;
                reg_next.bram_address <= (OTHERS => '0');
                reg_next.state <= wait_for_new_frame;

            WHEN OTHERS => NULL;
        END CASE;
    END PROCESS;

END ARCHITECTURE;